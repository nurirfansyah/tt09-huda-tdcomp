magic
tech sky130A
magscale 1 2
timestamp 1731262622
<< dnwell >>
rect -4234 -3709 9311 2246
<< nwell >>
rect 7237 -446 8275 129
rect -3854 -546 6074 -544
rect -3854 -840 6110 -546
rect -3818 -842 6110 -840
rect 6444 -1012 8275 -446
rect 7237 -2165 8275 -1012
<< locali >>
rect 6316 -434 6354 -400
rect 6388 -434 6426 -400
rect 6460 -434 6498 -400
rect 6532 -434 6570 -400
rect 6604 -434 6642 -400
rect 6676 -434 6714 -400
rect 6748 -434 6786 -400
rect 6316 -1058 6354 -1024
rect 6388 -1058 6426 -1024
rect 6460 -1058 6498 -1024
rect 6532 -1058 6570 -1024
rect 6604 -1058 6642 -1024
rect 6676 -1058 6714 -1024
rect 6748 -1058 6786 -1024
<< viali >>
rect 6282 -434 6316 -400
rect 6354 -434 6388 -400
rect 6426 -434 6460 -400
rect 6498 -434 6532 -400
rect 6570 -434 6604 -400
rect 6642 -434 6676 -400
rect 6714 -434 6748 -400
rect 6786 -434 6820 -400
rect 6909 -440 6943 -406
rect 6282 -1058 6316 -1024
rect 6354 -1058 6388 -1024
rect 6426 -1058 6460 -1024
rect 6498 -1058 6532 -1024
rect 6570 -1058 6604 -1024
rect 6642 -1058 6676 -1024
rect 6714 -1058 6748 -1024
rect 6786 -1058 6820 -1024
rect 6909 -1052 6943 -1018
<< metal1 >>
rect 6068 2134 9029 2246
rect -4241 2058 -4141 2072
rect -4241 2006 -4217 2058
rect -4165 2006 -4141 2058
rect -4241 1992 -4141 2006
rect -4524 1328 -4384 1330
rect -4524 1212 -4512 1328
rect -4396 1212 -4384 1328
rect -4524 1210 -4384 1212
rect -4514 -998 -4394 1210
rect -4231 -849 -4151 1992
rect 6872 -233 6972 2134
rect 5996 -400 6832 -394
rect 5996 -434 6282 -400
rect 6316 -434 6354 -400
rect 6388 -434 6426 -400
rect 6460 -434 6498 -400
rect 6532 -434 6570 -400
rect 6604 -434 6642 -400
rect 6676 -434 6714 -400
rect 6748 -434 6786 -400
rect 6820 -434 6832 -400
rect 5996 -440 6832 -434
rect 6887 -446 6900 -394
rect 6952 -446 6965 -394
rect -4045 -548 -3945 -534
rect -4045 -600 -4021 -548
rect -3969 -600 -3945 -548
rect -4045 -614 -3945 -600
rect -4241 -863 -4141 -849
rect -4241 -915 -4217 -863
rect -4165 -915 -4141 -863
rect -4241 -929 -4141 -915
rect -4524 -1012 -4384 -998
rect -4524 -1064 -4512 -1012
rect -4460 -1064 -4448 -1012
rect -4396 -1064 -4384 -1012
rect -4524 -1078 -4384 -1064
rect -4514 -2673 -4394 -1078
rect -4524 -2675 -4384 -2673
rect -4524 -2791 -4512 -2675
rect -4396 -2791 -4384 -2675
rect -4524 -2793 -4384 -2791
rect -4035 -3455 -3955 -614
rect -3866 -706 7341 -671
rect -3866 -758 -3860 -706
rect -3808 -758 -3796 -706
rect -3744 -758 -3732 -706
rect -3680 -758 -3668 -706
rect -3616 -758 -3604 -706
rect -3552 -758 -3540 -706
rect -3488 -758 -3476 -706
rect -3424 -758 -3412 -706
rect -3360 -758 -3348 -706
rect -3296 -758 -3284 -706
rect -3232 -758 -3220 -706
rect -3168 -758 -3156 -706
rect -3104 -758 -3092 -706
rect -3040 -758 -3028 -706
rect -2976 -758 -2964 -706
rect -2912 -758 -2900 -706
rect -2848 -758 -2836 -706
rect -2784 -758 -2772 -706
rect -2720 -758 -2708 -706
rect -2656 -758 -2644 -706
rect -2592 -758 -2580 -706
rect -2528 -758 -2516 -706
rect -2464 -758 -2452 -706
rect -2400 -758 -2388 -706
rect -2336 -758 -2324 -706
rect -2272 -758 -2260 -706
rect -2208 -758 -2196 -706
rect -2144 -758 -2132 -706
rect -2080 -758 -2068 -706
rect -2016 -758 -2004 -706
rect -1952 -758 -1940 -706
rect -1888 -758 -1876 -706
rect -1824 -758 -1812 -706
rect -1760 -758 -1748 -706
rect -1696 -758 -1684 -706
rect -1632 -758 -1620 -706
rect -1568 -758 -1556 -706
rect -1504 -758 -1492 -706
rect -1440 -758 -1428 -706
rect -1376 -758 -1364 -706
rect -1312 -758 -1300 -706
rect -1248 -758 -1236 -706
rect -1184 -758 -1172 -706
rect -1120 -758 -1108 -706
rect -1056 -758 -1044 -706
rect -992 -758 -980 -706
rect -928 -758 -916 -706
rect -864 -758 -852 -706
rect -800 -758 -788 -706
rect -736 -758 -724 -706
rect -672 -758 -660 -706
rect -608 -758 -596 -706
rect -544 -758 -532 -706
rect -480 -758 -468 -706
rect -416 -758 -404 -706
rect -352 -758 -340 -706
rect -288 -758 -276 -706
rect -224 -758 -212 -706
rect -160 -758 -148 -706
rect -96 -758 -84 -706
rect -32 -758 -20 -706
rect 32 -758 44 -706
rect 96 -758 108 -706
rect 160 -758 172 -706
rect 224 -758 236 -706
rect 288 -758 300 -706
rect 352 -758 364 -706
rect 416 -758 428 -706
rect 480 -758 492 -706
rect 544 -758 556 -706
rect 608 -758 620 -706
rect 672 -758 684 -706
rect 736 -758 748 -706
rect 800 -758 812 -706
rect 864 -758 876 -706
rect 928 -758 940 -706
rect 992 -758 1004 -706
rect 1056 -758 1068 -706
rect 1120 -758 1132 -706
rect 1184 -758 1196 -706
rect 1248 -758 1260 -706
rect 1312 -758 1324 -706
rect 1376 -758 1388 -706
rect 1440 -758 1452 -706
rect 1504 -758 1516 -706
rect 1568 -758 1580 -706
rect 1632 -758 1644 -706
rect 1696 -758 1708 -706
rect 1760 -758 1772 -706
rect 1824 -758 1836 -706
rect 1888 -758 1900 -706
rect 1952 -758 1964 -706
rect 2016 -758 2028 -706
rect 2080 -758 2092 -706
rect 2144 -758 2156 -706
rect 2208 -758 2220 -706
rect 2272 -758 2284 -706
rect 2336 -758 2348 -706
rect 2400 -758 2412 -706
rect 2464 -758 2476 -706
rect 2528 -758 2540 -706
rect 2592 -758 2604 -706
rect 2656 -758 2668 -706
rect 2720 -758 2732 -706
rect 2784 -758 2796 -706
rect 2848 -758 2860 -706
rect 2912 -758 2924 -706
rect 2976 -758 2988 -706
rect 3040 -758 3052 -706
rect 3104 -758 3116 -706
rect 3168 -758 3180 -706
rect 3232 -758 3244 -706
rect 3296 -758 3308 -706
rect 3360 -758 3372 -706
rect 3424 -758 3436 -706
rect 3488 -758 3500 -706
rect 3552 -758 3564 -706
rect 3616 -758 3628 -706
rect 3680 -758 3692 -706
rect 3744 -758 3756 -706
rect 3808 -758 3820 -706
rect 3872 -758 3884 -706
rect 3936 -758 3948 -706
rect 4000 -758 4012 -706
rect 4064 -758 4076 -706
rect 4128 -758 4140 -706
rect 4192 -758 4204 -706
rect 4256 -758 4268 -706
rect 4320 -758 4332 -706
rect 4384 -758 4396 -706
rect 4448 -758 4460 -706
rect 4512 -758 4524 -706
rect 4576 -758 4588 -706
rect 4640 -758 4652 -706
rect 4704 -758 4716 -706
rect 4768 -758 4780 -706
rect 4832 -758 4844 -706
rect 4896 -758 4908 -706
rect 4960 -758 4972 -706
rect 5024 -758 5036 -706
rect 5088 -758 5100 -706
rect 5152 -758 5164 -706
rect 5216 -758 5228 -706
rect 5280 -758 5292 -706
rect 5344 -758 5356 -706
rect 5408 -758 5420 -706
rect 5472 -758 5484 -706
rect 5536 -758 5548 -706
rect 5600 -758 5612 -706
rect 5664 -758 5676 -706
rect 5728 -758 5740 -706
rect 5792 -758 5804 -706
rect 5856 -758 5868 -706
rect 5920 -758 5932 -706
rect 5984 -758 5996 -706
rect 6048 -758 6060 -706
rect 6112 -758 6124 -706
rect 6176 -758 6188 -706
rect 6240 -758 6252 -706
rect 6304 -758 6316 -706
rect 6368 -758 6380 -706
rect 6432 -758 6444 -706
rect 6496 -758 6508 -706
rect 6560 -758 6572 -706
rect 6624 -758 6636 -706
rect 6688 -758 6700 -706
rect 6752 -758 6764 -706
rect 6816 -758 6828 -706
rect 6880 -758 6892 -706
rect 6944 -758 6956 -706
rect 7008 -758 7020 -706
rect 7072 -758 7084 -706
rect 7136 -758 7148 -706
rect 7200 -758 7212 -706
rect 7264 -758 7276 -706
rect 7328 -758 7341 -706
rect -3866 -791 7341 -758
rect 5935 -1024 6832 -1018
rect 5935 -1058 6282 -1024
rect 6316 -1058 6354 -1024
rect 6388 -1058 6426 -1024
rect 6460 -1058 6498 -1024
rect 6532 -1058 6570 -1024
rect 6604 -1058 6642 -1024
rect 6676 -1058 6714 -1024
rect 6748 -1058 6786 -1024
rect 6820 -1058 6832 -1024
rect 6887 -1058 6900 -1006
rect 6952 -1058 6965 -1006
rect 5935 -1064 6832 -1058
rect -4045 -3469 -3945 -3455
rect -4045 -3521 -4021 -3469
rect -3969 -3521 -3945 -3469
rect -4045 -3535 -3945 -3521
rect 6871 -3597 6971 -1225
rect 8932 -3597 9029 2134
rect 6115 -3709 9029 -3597
<< via1 >>
rect -4217 2006 -4165 2058
rect -4512 1212 -4396 1328
rect 6900 -406 6952 -394
rect 6900 -440 6909 -406
rect 6909 -440 6943 -406
rect 6943 -440 6952 -406
rect 6900 -446 6952 -440
rect -4021 -600 -3969 -548
rect -4217 -915 -4165 -863
rect -4512 -1064 -4460 -1012
rect -4448 -1064 -4396 -1012
rect -4512 -2791 -4396 -2675
rect -3860 -758 -3808 -706
rect -3796 -758 -3744 -706
rect -3732 -758 -3680 -706
rect -3668 -758 -3616 -706
rect -3604 -758 -3552 -706
rect -3540 -758 -3488 -706
rect -3476 -758 -3424 -706
rect -3412 -758 -3360 -706
rect -3348 -758 -3296 -706
rect -3284 -758 -3232 -706
rect -3220 -758 -3168 -706
rect -3156 -758 -3104 -706
rect -3092 -758 -3040 -706
rect -3028 -758 -2976 -706
rect -2964 -758 -2912 -706
rect -2900 -758 -2848 -706
rect -2836 -758 -2784 -706
rect -2772 -758 -2720 -706
rect -2708 -758 -2656 -706
rect -2644 -758 -2592 -706
rect -2580 -758 -2528 -706
rect -2516 -758 -2464 -706
rect -2452 -758 -2400 -706
rect -2388 -758 -2336 -706
rect -2324 -758 -2272 -706
rect -2260 -758 -2208 -706
rect -2196 -758 -2144 -706
rect -2132 -758 -2080 -706
rect -2068 -758 -2016 -706
rect -2004 -758 -1952 -706
rect -1940 -758 -1888 -706
rect -1876 -758 -1824 -706
rect -1812 -758 -1760 -706
rect -1748 -758 -1696 -706
rect -1684 -758 -1632 -706
rect -1620 -758 -1568 -706
rect -1556 -758 -1504 -706
rect -1492 -758 -1440 -706
rect -1428 -758 -1376 -706
rect -1364 -758 -1312 -706
rect -1300 -758 -1248 -706
rect -1236 -758 -1184 -706
rect -1172 -758 -1120 -706
rect -1108 -758 -1056 -706
rect -1044 -758 -992 -706
rect -980 -758 -928 -706
rect -916 -758 -864 -706
rect -852 -758 -800 -706
rect -788 -758 -736 -706
rect -724 -758 -672 -706
rect -660 -758 -608 -706
rect -596 -758 -544 -706
rect -532 -758 -480 -706
rect -468 -758 -416 -706
rect -404 -758 -352 -706
rect -340 -758 -288 -706
rect -276 -758 -224 -706
rect -212 -758 -160 -706
rect -148 -758 -96 -706
rect -84 -758 -32 -706
rect -20 -758 32 -706
rect 44 -758 96 -706
rect 108 -758 160 -706
rect 172 -758 224 -706
rect 236 -758 288 -706
rect 300 -758 352 -706
rect 364 -758 416 -706
rect 428 -758 480 -706
rect 492 -758 544 -706
rect 556 -758 608 -706
rect 620 -758 672 -706
rect 684 -758 736 -706
rect 748 -758 800 -706
rect 812 -758 864 -706
rect 876 -758 928 -706
rect 940 -758 992 -706
rect 1004 -758 1056 -706
rect 1068 -758 1120 -706
rect 1132 -758 1184 -706
rect 1196 -758 1248 -706
rect 1260 -758 1312 -706
rect 1324 -758 1376 -706
rect 1388 -758 1440 -706
rect 1452 -758 1504 -706
rect 1516 -758 1568 -706
rect 1580 -758 1632 -706
rect 1644 -758 1696 -706
rect 1708 -758 1760 -706
rect 1772 -758 1824 -706
rect 1836 -758 1888 -706
rect 1900 -758 1952 -706
rect 1964 -758 2016 -706
rect 2028 -758 2080 -706
rect 2092 -758 2144 -706
rect 2156 -758 2208 -706
rect 2220 -758 2272 -706
rect 2284 -758 2336 -706
rect 2348 -758 2400 -706
rect 2412 -758 2464 -706
rect 2476 -758 2528 -706
rect 2540 -758 2592 -706
rect 2604 -758 2656 -706
rect 2668 -758 2720 -706
rect 2732 -758 2784 -706
rect 2796 -758 2848 -706
rect 2860 -758 2912 -706
rect 2924 -758 2976 -706
rect 2988 -758 3040 -706
rect 3052 -758 3104 -706
rect 3116 -758 3168 -706
rect 3180 -758 3232 -706
rect 3244 -758 3296 -706
rect 3308 -758 3360 -706
rect 3372 -758 3424 -706
rect 3436 -758 3488 -706
rect 3500 -758 3552 -706
rect 3564 -758 3616 -706
rect 3628 -758 3680 -706
rect 3692 -758 3744 -706
rect 3756 -758 3808 -706
rect 3820 -758 3872 -706
rect 3884 -758 3936 -706
rect 3948 -758 4000 -706
rect 4012 -758 4064 -706
rect 4076 -758 4128 -706
rect 4140 -758 4192 -706
rect 4204 -758 4256 -706
rect 4268 -758 4320 -706
rect 4332 -758 4384 -706
rect 4396 -758 4448 -706
rect 4460 -758 4512 -706
rect 4524 -758 4576 -706
rect 4588 -758 4640 -706
rect 4652 -758 4704 -706
rect 4716 -758 4768 -706
rect 4780 -758 4832 -706
rect 4844 -758 4896 -706
rect 4908 -758 4960 -706
rect 4972 -758 5024 -706
rect 5036 -758 5088 -706
rect 5100 -758 5152 -706
rect 5164 -758 5216 -706
rect 5228 -758 5280 -706
rect 5292 -758 5344 -706
rect 5356 -758 5408 -706
rect 5420 -758 5472 -706
rect 5484 -758 5536 -706
rect 5548 -758 5600 -706
rect 5612 -758 5664 -706
rect 5676 -758 5728 -706
rect 5740 -758 5792 -706
rect 5804 -758 5856 -706
rect 5868 -758 5920 -706
rect 5932 -758 5984 -706
rect 5996 -758 6048 -706
rect 6060 -758 6112 -706
rect 6124 -758 6176 -706
rect 6188 -758 6240 -706
rect 6252 -758 6304 -706
rect 6316 -758 6368 -706
rect 6380 -758 6432 -706
rect 6444 -758 6496 -706
rect 6508 -758 6560 -706
rect 6572 -758 6624 -706
rect 6636 -758 6688 -706
rect 6700 -758 6752 -706
rect 6764 -758 6816 -706
rect 6828 -758 6880 -706
rect 6892 -758 6944 -706
rect 6956 -758 7008 -706
rect 7020 -758 7072 -706
rect 7084 -758 7136 -706
rect 7148 -758 7200 -706
rect 7212 -758 7264 -706
rect 7276 -758 7328 -706
rect 6900 -1018 6952 -1006
rect 6900 -1052 6909 -1018
rect 6909 -1052 6943 -1018
rect 6943 -1052 6952 -1018
rect 6900 -1058 6952 -1052
rect -4021 -3521 -3969 -3469
<< metal2 >>
rect -4231 2072 -4151 2082
rect -4231 2058 -3775 2072
rect -4231 2006 -4217 2058
rect -4165 2006 -3775 2058
rect -4231 1992 -3775 2006
rect -4231 1982 -4151 1992
rect -4514 1330 -4394 1340
rect -4514 1328 -3735 1330
rect -4514 1212 -4512 1328
rect -4396 1212 -3735 1328
rect -4514 1210 -3735 1212
rect -4514 1200 -4394 1210
rect 8422 -216 9311 -164
rect 8422 -247 8474 -216
rect 6897 -394 6955 -384
rect 6897 -446 6900 -394
rect 6952 -395 6955 -394
rect 7420 -393 7476 -383
rect 6952 -446 7420 -395
rect 6897 -456 6955 -446
rect 7476 -446 7492 -395
rect 7420 -459 7476 -449
rect -4035 -534 -3955 -524
rect -4836 -548 -3774 -534
rect -4836 -600 -4021 -548
rect -3969 -600 -3774 -548
rect -4836 -614 -3774 -600
rect -4035 -624 -3955 -614
rect -3987 -684 7340 -676
rect -4836 -706 7340 -684
rect -4836 -758 -3860 -706
rect -3808 -758 -3796 -706
rect -3744 -758 -3732 -706
rect -3680 -758 -3668 -706
rect -3616 -758 -3604 -706
rect -3552 -758 -3540 -706
rect -3488 -758 -3476 -706
rect -3424 -758 -3412 -706
rect -3360 -758 -3348 -706
rect -3296 -758 -3284 -706
rect -3232 -758 -3220 -706
rect -3168 -758 -3156 -706
rect -3104 -758 -3092 -706
rect -3040 -758 -3028 -706
rect -2976 -758 -2964 -706
rect -2912 -758 -2900 -706
rect -2848 -758 -2836 -706
rect -2784 -758 -2772 -706
rect -2720 -758 -2708 -706
rect -2656 -758 -2644 -706
rect -2592 -758 -2580 -706
rect -2528 -758 -2516 -706
rect -2464 -758 -2452 -706
rect -2400 -758 -2388 -706
rect -2336 -758 -2324 -706
rect -2272 -758 -2260 -706
rect -2208 -758 -2196 -706
rect -2144 -758 -2132 -706
rect -2080 -758 -2068 -706
rect -2016 -758 -2004 -706
rect -1952 -758 -1940 -706
rect -1888 -758 -1876 -706
rect -1824 -758 -1812 -706
rect -1760 -758 -1748 -706
rect -1696 -758 -1684 -706
rect -1632 -758 -1620 -706
rect -1568 -758 -1556 -706
rect -1504 -758 -1492 -706
rect -1440 -758 -1428 -706
rect -1376 -758 -1364 -706
rect -1312 -758 -1300 -706
rect -1248 -758 -1236 -706
rect -1184 -758 -1172 -706
rect -1120 -758 -1108 -706
rect -1056 -758 -1044 -706
rect -992 -758 -980 -706
rect -928 -758 -916 -706
rect -864 -758 -852 -706
rect -800 -758 -788 -706
rect -736 -758 -724 -706
rect -672 -758 -660 -706
rect -608 -758 -596 -706
rect -544 -758 -532 -706
rect -480 -758 -468 -706
rect -416 -758 -404 -706
rect -352 -758 -340 -706
rect -288 -758 -276 -706
rect -224 -758 -212 -706
rect -160 -758 -148 -706
rect -96 -758 -84 -706
rect -32 -758 -20 -706
rect 32 -758 44 -706
rect 96 -758 108 -706
rect 160 -758 172 -706
rect 224 -758 236 -706
rect 288 -758 300 -706
rect 352 -758 364 -706
rect 416 -758 428 -706
rect 480 -758 492 -706
rect 544 -758 556 -706
rect 608 -758 620 -706
rect 672 -758 684 -706
rect 736 -758 748 -706
rect 800 -758 812 -706
rect 864 -758 876 -706
rect 928 -758 940 -706
rect 992 -758 1004 -706
rect 1056 -758 1068 -706
rect 1120 -758 1132 -706
rect 1184 -758 1196 -706
rect 1248 -758 1260 -706
rect 1312 -758 1324 -706
rect 1376 -758 1388 -706
rect 1440 -758 1452 -706
rect 1504 -758 1516 -706
rect 1568 -758 1580 -706
rect 1632 -758 1644 -706
rect 1696 -758 1708 -706
rect 1760 -758 1772 -706
rect 1824 -758 1836 -706
rect 1888 -758 1900 -706
rect 1952 -758 1964 -706
rect 2016 -758 2028 -706
rect 2080 -758 2092 -706
rect 2144 -758 2156 -706
rect 2208 -758 2220 -706
rect 2272 -758 2284 -706
rect 2336 -758 2348 -706
rect 2400 -758 2412 -706
rect 2464 -758 2476 -706
rect 2528 -758 2540 -706
rect 2592 -758 2604 -706
rect 2656 -758 2668 -706
rect 2720 -758 2732 -706
rect 2784 -758 2796 -706
rect 2848 -758 2860 -706
rect 2912 -758 2924 -706
rect 2976 -758 2988 -706
rect 3040 -758 3052 -706
rect 3104 -758 3116 -706
rect 3168 -758 3180 -706
rect 3232 -758 3244 -706
rect 3296 -758 3308 -706
rect 3360 -758 3372 -706
rect 3424 -758 3436 -706
rect 3488 -758 3500 -706
rect 3552 -758 3564 -706
rect 3616 -758 3628 -706
rect 3680 -758 3692 -706
rect 3744 -758 3756 -706
rect 3808 -758 3820 -706
rect 3872 -758 3884 -706
rect 3936 -758 3948 -706
rect 4000 -758 4012 -706
rect 4064 -758 4076 -706
rect 4128 -758 4140 -706
rect 4192 -758 4204 -706
rect 4256 -758 4268 -706
rect 4320 -758 4332 -706
rect 4384 -758 4396 -706
rect 4448 -758 4460 -706
rect 4512 -758 4524 -706
rect 4576 -758 4588 -706
rect 4640 -758 4652 -706
rect 4704 -758 4716 -706
rect 4768 -758 4780 -706
rect 4832 -758 4844 -706
rect 4896 -758 4908 -706
rect 4960 -758 4972 -706
rect 5024 -758 5036 -706
rect 5088 -758 5100 -706
rect 5152 -758 5164 -706
rect 5216 -758 5228 -706
rect 5280 -758 5292 -706
rect 5344 -758 5356 -706
rect 5408 -758 5420 -706
rect 5472 -758 5484 -706
rect 5536 -758 5548 -706
rect 5600 -758 5612 -706
rect 5664 -758 5676 -706
rect 5728 -758 5740 -706
rect 5792 -758 5804 -706
rect 5856 -758 5868 -706
rect 5920 -758 5932 -706
rect 5984 -758 5996 -706
rect 6048 -758 6060 -706
rect 6112 -758 6124 -706
rect 6176 -758 6188 -706
rect 6240 -758 6252 -706
rect 6304 -758 6316 -706
rect 6368 -758 6380 -706
rect 6432 -758 6444 -706
rect 6496 -758 6508 -706
rect 6560 -758 6572 -706
rect 6624 -758 6636 -706
rect 6688 -758 6700 -706
rect 6752 -758 6764 -706
rect 6816 -758 6828 -706
rect 6880 -758 6892 -706
rect 6944 -758 6956 -706
rect 7008 -758 7020 -706
rect 7072 -758 7084 -706
rect 7136 -758 7148 -706
rect 7200 -758 7212 -706
rect 7264 -758 7276 -706
rect 7328 -758 7340 -706
rect -4836 -779 7340 -758
rect -3987 -788 7340 -779
rect -4231 -849 -4151 -839
rect -4836 -863 -3774 -849
rect -4836 -915 -4217 -863
rect -4165 -915 -3774 -863
rect -4836 -929 -3774 -915
rect -4231 -939 -4151 -929
rect -4514 -998 -4394 -988
rect -4836 -1012 -4394 -998
rect -4836 -1064 -4512 -1012
rect -4460 -1064 -4448 -1012
rect -4396 -1064 -4394 -1012
rect -4836 -1078 -4394 -1064
rect 6897 -1006 6955 -996
rect 6897 -1058 6900 -1006
rect 6952 -1058 7619 -1006
rect 6897 -1068 6955 -1058
rect -4514 -1088 -4394 -1078
rect 8427 -1241 8483 -1203
rect 8427 -1297 9311 -1241
rect -4514 -2673 -4394 -2663
rect -4514 -2675 -3735 -2673
rect -4514 -2791 -4512 -2675
rect -4396 -2791 -3735 -2675
rect -4514 -2793 -3735 -2791
rect -4514 -2803 -4394 -2793
rect -4035 -3455 -3955 -3445
rect -4035 -3469 -3775 -3455
rect -4035 -3521 -4021 -3469
rect -3969 -3521 -3775 -3469
rect -4035 -3535 -3775 -3521
rect -4035 -3545 -3955 -3535
<< via2 >>
rect 7420 -449 7476 -393
<< metal3 >>
rect 7410 -393 7486 -318
rect 7410 -449 7420 -393
rect 7476 -449 7486 -393
rect 7410 -454 7486 -449
use delay_element  delay_element_0
timestamp 1731262622
transform 1 0 -3748 0 1 -1956
box -119 -1753 9905 1280
use delay_element  delay_element_1
timestamp 1731262622
transform 1 0 -3748 0 -1 493
box -119 -1753 9905 1280
use phase_detector  phase_detector_0
timestamp 1731262622
transform 0 -1 9209 -1 0 -453
box -1184 180 1722 1972
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1731262622
transform -1 0 6972 0 1 -1273
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_1
timestamp 1731262622
transform -1 0 6972 0 -1 -185
box -38 -48 866 592
<< labels >>
flabel metal2 s 9256 -207 9301 -173 0 FreeSans 1250 0 0 0 outp
port 1 nsew
flabel metal2 s 9254 -1285 9299 -1251 0 FreeSans 1250 0 0 0 outn
port 2 nsew
flabel metal2 s -3831 -747 -3786 -713 0 FreeSans 1250 0 0 0 vdda
port 3 nsew
flabel metal2 s -4807 -1058 -4762 -1024 0 FreeSans 1250 0 0 0 start
port 4 nsew
flabel metal2 s -4808 -598 -4766 -546 0 FreeSans 1250 0 0 0 vinn
port 5 nsew
flabel metal2 s -4816 -914 -4758 -860 0 FreeSans 1250 0 0 0 vinp
port 6 nsew
flabel metal1 s 6878 -3686 6962 -3612 0 FreeSans 1250 0 0 0 vssa
port 7 nsew
<< end >>
