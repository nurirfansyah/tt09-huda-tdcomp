magic
tech sky130A
magscale 1 2
timestamp 1731261117
<< dnwell >>
rect -4234 -3709 9311 2246
<< nwell >>
rect 7237 -446 8275 129
rect -3854 -546 6074 -544
rect -3854 -840 6110 -546
rect -3818 -842 6110 -840
rect 6444 -1012 8275 -446
rect 7237 -2165 8275 -1012
<< viali >>
rect 6282 -434 6820 -400
rect 6909 -440 6943 -406
rect 6282 -1058 6820 -1024
rect 6909 -1052 6943 -1018
<< metal1 >>
rect 6068 2134 9029 2246
rect -4241 1992 -4231 2072
rect -4151 1992 -4141 2072
rect -4524 1210 -4514 1330
rect -4394 1210 -4384 1330
rect -4514 -998 -4394 1210
rect -4231 -849 -4151 1992
rect 6872 -233 6972 2134
rect 5996 -400 6832 -394
rect 5996 -434 6282 -400
rect 6820 -434 6832 -400
rect 5996 -440 6832 -434
rect 6887 -446 6897 -394
rect 6955 -446 6965 -394
rect -4045 -614 -4035 -534
rect -3955 -614 -3945 -534
rect -4241 -929 -4231 -849
rect -4151 -929 -4141 -849
rect -4524 -1078 -4514 -998
rect -4394 -1078 -4384 -998
rect -4514 -2673 -4394 -1078
rect -4524 -2793 -4514 -2673
rect -4394 -2793 -4384 -2673
rect -4035 -3455 -3955 -614
rect -3866 -684 7341 -671
rect 7334 -779 7341 -684
rect -3866 -791 7341 -779
rect 5935 -1024 6832 -1018
rect 5935 -1058 6282 -1024
rect 6820 -1058 6832 -1024
rect 6887 -1058 6897 -1006
rect 6955 -1058 6965 -1006
rect 5935 -1064 6832 -1058
rect -4045 -3535 -4035 -3455
rect -3955 -3535 -3945 -3455
rect 6871 -3597 6971 -1225
rect 8932 -3597 9029 2134
rect 6115 -3709 9029 -3597
<< via1 >>
rect -4231 1992 -4151 2072
rect -4514 1210 -4394 1330
rect 6897 -406 6955 -394
rect 6897 -440 6909 -406
rect 6909 -440 6943 -406
rect 6943 -440 6955 -406
rect 6897 -446 6955 -440
rect -4035 -614 -3955 -534
rect -4231 -929 -4151 -849
rect -4514 -1078 -4394 -998
rect -4514 -2793 -4394 -2673
rect -3866 -779 7334 -684
rect 6897 -1018 6955 -1006
rect 6897 -1052 6909 -1018
rect 6909 -1052 6943 -1018
rect 6943 -1052 6955 -1018
rect 6897 -1058 6955 -1052
rect -4035 -3535 -3955 -3455
<< metal2 >>
rect -4231 2072 -4151 2082
rect -4151 1992 -3775 2072
rect -4231 1982 -4151 1992
rect -4514 1330 -4394 1340
rect -4394 1210 -3735 1330
rect -4514 1200 -4394 1210
rect 8422 -216 9311 -164
rect 8422 -247 8474 -216
rect 6897 -394 6955 -384
rect 7420 -393 7476 -383
rect 6955 -446 7420 -395
rect 6897 -456 6955 -446
rect 7476 -446 7492 -395
rect 7420 -459 7476 -449
rect -4035 -534 -3955 -524
rect -4836 -614 -4035 -534
rect -3955 -614 -3774 -534
rect -4035 -624 -3955 -614
rect -3987 -684 7340 -676
rect -4836 -779 -3866 -684
rect 7334 -779 7340 -684
rect -3987 -788 7340 -779
rect -4231 -849 -4151 -839
rect -4836 -929 -4231 -849
rect -4151 -929 -3774 -849
rect -4231 -939 -4151 -929
rect -4514 -998 -4394 -988
rect -4836 -1078 -4514 -998
rect 6897 -1006 6955 -996
rect 6955 -1058 7619 -1006
rect 6897 -1068 6955 -1058
rect -4514 -1088 -4394 -1078
rect 8427 -1241 8483 -1203
rect 8427 -1297 9311 -1241
rect -4514 -2673 -4394 -2663
rect -4394 -2793 -3735 -2673
rect -4514 -2803 -4394 -2793
rect -4035 -3455 -3955 -3445
rect -3955 -3535 -3775 -3455
rect -4035 -3545 -3955 -3535
<< via2 >>
rect 7420 -449 7476 -393
<< metal3 >>
rect 7410 -393 7486 -318
rect 7410 -449 7420 -393
rect 7476 -449 7486 -393
rect 7410 -454 7486 -449
use delay_element  delay_element_0
timestamp 1731173062
transform 1 0 -3748 0 1 -1956
box -119 -1753 9905 1280
use delay_element  delay_element_1
timestamp 1731173062
transform 1 0 -3748 0 -1 493
box -119 -1753 9905 1280
use phase_detector  phase_detector_0
timestamp 1731258661
transform 0 -1 9209 -1 0 -453
box -1184 180 1722 1972
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform -1 0 6972 0 1 -1273
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_1
timestamp 1730246015
transform -1 0 6972 0 -1 -185
box -38 -48 866 592
<< labels >>
flabel metal2 9256 -207 9301 -173 0 FreeSans 800 0 0 0 outp
port 0 nsew
flabel metal2 9254 -1285 9299 -1251 0 FreeSans 800 0 0 0 outn
port 1 nsew
flabel metal2 -4807 -1058 -4762 -1024 0 FreeSans 800 0 0 0 start
port 5 nsew
flabel metal2 -4808 -598 -4766 -546 0 FreeSans 800 0 0 0 vinn
port 9 nsew
flabel metal2 -4816 -914 -4758 -860 0 FreeSans 800 0 0 0 vinp
port 11 nsew
flabel metal1 6878 -3686 6962 -3612 0 FreeSans 800 0 0 0 vssa
port 13 nsew
flabel via1 -3831 -747 -3786 -713 0 FreeSans 800 0 0 0 vdda
port 2 nsew
<< end >>
