magic
tech sky130A
magscale 1 2
timestamp 1731262622
<< nwell >>
rect -1174 918 1367 1956
rect 199 905 372 918
<< locali >>
rect -1042 1902 -1032 1936
rect -998 1902 -960 1936
rect -926 1902 -888 1936
rect -854 1902 -816 1936
rect -782 1902 -744 1936
rect -710 1902 -672 1936
rect -638 1902 -600 1936
rect -566 1902 -528 1936
rect -494 1902 -456 1936
rect -422 1902 -384 1936
rect -350 1902 -312 1936
rect -278 1902 -268 1936
rect 806 1902 816 1936
rect 850 1902 888 1936
rect 922 1902 960 1936
rect 994 1902 1032 1936
rect 1066 1902 1104 1936
rect 1138 1902 1176 1936
rect 1210 1902 1248 1936
rect 1282 1902 1320 1936
rect 1354 1902 1392 1936
rect 1426 1902 1464 1936
rect 1498 1902 1536 1936
rect 1570 1902 1580 1936
rect -1042 216 -1025 250
rect -991 216 -953 250
rect -919 216 -881 250
rect -847 216 -809 250
rect -775 216 -737 250
rect -703 216 -686 250
rect 1224 216 1241 250
rect 1275 216 1313 250
rect 1347 216 1385 250
rect 1419 216 1457 250
rect 1491 216 1529 250
rect 1563 216 1580 250
<< viali >>
rect -1032 1902 -998 1936
rect -960 1902 -926 1936
rect -888 1902 -854 1936
rect -816 1902 -782 1936
rect -744 1902 -710 1936
rect -672 1902 -638 1936
rect -600 1902 -566 1936
rect -528 1902 -494 1936
rect -456 1902 -422 1936
rect -384 1902 -350 1936
rect -312 1902 -278 1936
rect 816 1902 850 1936
rect 888 1902 922 1936
rect 960 1902 994 1936
rect 1032 1902 1066 1936
rect 1104 1902 1138 1936
rect 1176 1902 1210 1936
rect 1248 1902 1282 1936
rect 1320 1902 1354 1936
rect 1392 1902 1426 1936
rect 1464 1902 1498 1936
rect 1536 1902 1570 1936
rect 483 1027 517 1061
rect -62 859 -28 893
rect 106 859 140 893
rect 396 859 430 893
rect 564 859 598 893
rect 109 737 143 771
rect 525 737 559 771
rect -1025 216 -991 250
rect -953 216 -919 250
rect -881 216 -847 250
rect -809 216 -775 250
rect -737 216 -703 250
rect 1241 216 1275 250
rect 1313 216 1347 250
rect 1385 216 1419 250
rect 1457 216 1491 250
rect 1529 216 1563 250
<< metal1 >>
rect -1174 1936 1712 1972
rect -1174 1902 -1032 1936
rect -998 1902 -960 1936
rect -926 1902 -888 1936
rect -854 1902 -816 1936
rect -782 1902 -744 1936
rect -710 1902 -672 1936
rect -638 1902 -600 1936
rect -566 1902 -528 1936
rect -494 1902 -456 1936
rect -422 1902 -384 1936
rect -350 1902 -312 1936
rect -278 1902 816 1936
rect 850 1902 888 1936
rect 922 1902 960 1936
rect 994 1902 1032 1936
rect 1066 1902 1104 1936
rect 1138 1902 1176 1936
rect 1210 1902 1248 1936
rect 1282 1902 1320 1936
rect 1354 1902 1392 1936
rect 1426 1902 1464 1936
rect 1498 1902 1536 1936
rect 1570 1902 1712 1936
rect -1174 1875 1712 1902
rect -1062 1787 -986 1794
rect -1062 1735 -1050 1787
rect -998 1735 -986 1787
rect -405 1782 -355 1875
rect -324 1787 -248 1794
rect -1062 1728 -986 1735
rect -1184 1471 -1108 1478
rect -1184 1419 -1172 1471
rect -1120 1419 -1108 1471
rect -1184 1412 -1108 1419
rect -1062 1471 -986 1478
rect -1062 1419 -1050 1471
rect -998 1419 -986 1471
rect -955 1466 -905 1740
rect -324 1735 -312 1787
rect -260 1735 -248 1787
rect -324 1728 -248 1735
rect -314 1656 -258 1728
rect -324 1649 -248 1656
rect -324 1597 -312 1649
rect -260 1597 -248 1649
rect -324 1590 -248 1597
rect -324 1471 -248 1478
rect -1062 1412 -986 1419
rect -1174 424 -1122 1412
rect -407 1322 -355 1425
rect -324 1419 -312 1471
rect -260 1419 -248 1471
rect -324 1412 -248 1419
rect -417 1270 -407 1322
rect -355 1270 -345 1322
rect -208 1270 -198 1322
rect -146 1270 -136 1322
rect -1052 882 -996 1162
rect -417 1150 -407 1202
rect -355 1150 -345 1202
rect -814 1006 -764 1108
rect -314 1096 -258 1162
rect -198 1006 -146 1270
rect 573 1236 636 1875
rect 786 1787 862 1794
rect 786 1735 798 1787
rect 850 1735 862 1787
rect 893 1782 943 1875
rect 786 1728 862 1735
rect 674 1656 730 1666
rect 674 1649 754 1656
rect 674 1597 689 1649
rect 741 1597 754 1649
rect 674 1590 754 1597
rect 674 1478 730 1590
rect 664 1471 740 1478
rect 664 1419 676 1471
rect 728 1419 740 1471
rect 664 1412 740 1419
rect 786 1471 862 1478
rect 786 1419 798 1471
rect 850 1419 862 1471
rect 1443 1466 1493 1740
rect 1534 1728 1590 1794
rect 1524 1471 1600 1478
rect 786 1412 862 1419
rect 893 1322 945 1424
rect 1524 1419 1536 1471
rect 1588 1419 1600 1471
rect 1524 1412 1600 1419
rect 1646 1471 1722 1478
rect 1646 1419 1658 1471
rect 1710 1419 1722 1471
rect 1646 1412 1722 1419
rect 674 1270 684 1322
rect 736 1270 746 1322
rect 883 1270 893 1322
rect 945 1270 955 1322
rect -98 1184 -72 1236
rect -20 1184 113 1236
rect 165 1184 389 1236
rect 441 1184 573 1236
rect 625 1184 636 1236
rect -98 1140 636 1184
rect 461 1098 539 1100
rect 461 1077 474 1098
rect 90 1046 474 1077
rect 526 1046 539 1098
rect 90 1027 483 1046
rect 517 1044 539 1046
rect 517 1027 529 1044
rect 90 1010 529 1027
rect -824 954 -812 1006
rect -760 954 -748 1006
rect -208 954 -198 1006
rect -146 954 -136 1006
rect -91 975 -4 976
rect -1062 830 -1050 882
rect -998 830 -986 882
rect -1052 674 -996 830
rect -814 728 -764 954
rect -91 923 -74 975
rect -22 923 -4 975
rect -91 922 -4 923
rect -81 893 -14 922
rect -81 859 -62 893
rect -28 859 -14 893
rect -81 853 -14 859
rect 90 893 157 1010
rect 90 859 106 893
rect 140 859 157 893
rect 90 843 157 859
rect 238 893 446 904
rect 238 859 396 893
rect 430 859 446 893
rect 238 848 446 859
rect 538 902 625 909
rect 538 850 555 902
rect 607 850 625 902
rect 684 882 736 1270
rect 796 1096 852 1162
rect 883 1150 893 1202
rect 945 1150 955 1202
rect 1302 882 1352 1108
rect 1534 1006 1590 1162
rect 1524 954 1536 1006
rect 1588 954 1600 1006
rect 238 787 294 848
rect 538 843 625 850
rect 674 830 684 882
rect 736 830 746 882
rect 1286 830 1298 882
rect 1350 830 1362 882
rect 87 785 294 787
rect -1184 417 -1108 424
rect -1184 365 -1172 417
rect -1120 365 -1108 417
rect -1184 358 -1108 365
rect -1072 417 -996 424
rect -1072 365 -1060 417
rect -1008 365 -996 417
rect -814 412 -764 686
rect -732 674 -676 740
rect 87 733 100 785
rect 152 733 294 785
rect 87 731 294 733
rect 503 780 581 782
rect 503 728 516 780
rect 568 728 581 780
rect 503 726 581 728
rect -98 596 637 692
rect 1214 674 1270 740
rect 1302 728 1352 830
rect -1072 358 -996 365
rect -814 277 -764 370
rect -732 358 -676 424
rect 573 277 636 596
rect 1214 358 1270 424
rect 1302 412 1352 686
rect 1534 674 1590 954
rect 1660 424 1712 1412
rect 1534 417 1610 424
rect 1302 277 1352 368
rect 1534 365 1546 417
rect 1598 365 1610 417
rect 1534 358 1610 365
rect 1646 417 1722 424
rect 1646 365 1658 417
rect 1710 365 1722 417
rect 1646 358 1722 365
rect -1174 250 1712 277
rect -1174 216 -1025 250
rect -991 216 -953 250
rect -919 216 -881 250
rect -847 216 -809 250
rect -775 216 -737 250
rect -703 216 1241 250
rect 1275 216 1313 250
rect 1347 216 1385 250
rect 1419 216 1457 250
rect 1491 216 1529 250
rect 1563 216 1712 250
rect -1174 180 1712 216
<< via1 >>
rect -1050 1735 -998 1787
rect -1172 1419 -1120 1471
rect -1050 1419 -998 1471
rect -312 1735 -260 1787
rect -312 1597 -260 1649
rect -312 1419 -260 1471
rect -407 1270 -355 1322
rect -198 1270 -146 1322
rect -407 1150 -355 1202
rect 798 1735 850 1787
rect 689 1597 741 1649
rect 676 1419 728 1471
rect 798 1419 850 1471
rect 1536 1419 1588 1471
rect 1658 1419 1710 1471
rect 684 1270 736 1322
rect 893 1270 945 1322
rect -72 1184 -20 1236
rect 113 1184 165 1236
rect 389 1184 441 1236
rect 573 1184 625 1236
rect 474 1061 526 1098
rect 474 1046 483 1061
rect 483 1046 517 1061
rect 517 1046 526 1061
rect -812 954 -760 1006
rect -198 954 -146 1006
rect -1050 830 -998 882
rect -74 923 -22 975
rect 555 893 607 902
rect 555 859 564 893
rect 564 859 598 893
rect 598 859 607 893
rect 555 850 607 859
rect 893 1150 945 1202
rect 1536 954 1588 1006
rect 684 830 736 882
rect 1298 830 1350 882
rect -1172 365 -1120 417
rect -1060 365 -1008 417
rect 100 771 152 785
rect 100 737 109 771
rect 109 737 143 771
rect 143 737 152 771
rect 100 733 152 737
rect 516 771 568 780
rect 516 737 525 771
rect 525 737 559 771
rect 559 737 568 771
rect 516 728 568 737
rect 1546 365 1598 417
rect 1658 365 1710 417
<< metal2 >>
rect -1052 1794 -996 1804
rect -1174 1787 -996 1794
rect -1174 1735 -1050 1787
rect -998 1735 -996 1787
rect -1174 1728 -996 1735
rect -1052 1718 -996 1728
rect -314 1787 -258 1804
rect -314 1735 -312 1787
rect -260 1735 -258 1787
rect -314 1718 -258 1735
rect 796 1789 852 1804
rect 796 1718 852 1733
rect -314 1656 -258 1666
rect 687 1656 744 1666
rect -314 1649 744 1656
rect -314 1597 -312 1649
rect -260 1597 689 1649
rect 741 1597 744 1649
rect -314 1590 744 1597
rect -314 1580 -258 1590
rect 687 1580 744 1590
rect -1174 1478 -1118 1488
rect -1052 1478 -996 1488
rect -1174 1471 -996 1478
rect -1174 1419 -1172 1471
rect -1120 1419 -1050 1471
rect -998 1419 -996 1471
rect -1174 1412 -996 1419
rect -1174 1402 -1118 1412
rect -1052 1402 -996 1412
rect -314 1478 -258 1488
rect -192 1478 -136 1488
rect -314 1473 -136 1478
rect -314 1471 -192 1473
rect -314 1419 -312 1471
rect -260 1419 -192 1471
rect -314 1417 -192 1419
rect -314 1412 -136 1417
rect -314 1402 -258 1412
rect -192 1402 -136 1412
rect 674 1478 730 1488
rect 796 1478 852 1488
rect 674 1471 852 1478
rect 674 1419 676 1471
rect 728 1419 798 1471
rect 850 1419 852 1471
rect 674 1412 852 1419
rect 674 1402 730 1412
rect 796 1402 852 1412
rect 1534 1478 1590 1488
rect 1656 1478 1712 1488
rect 1534 1471 1712 1478
rect 1534 1419 1536 1471
rect 1588 1419 1658 1471
rect 1710 1419 1712 1471
rect 1534 1412 1712 1419
rect 1534 1402 1590 1412
rect 1656 1402 1712 1412
rect -407 1322 -355 1332
rect -198 1322 -146 1332
rect -355 1270 -198 1322
rect -407 1260 -355 1270
rect -198 1260 -146 1270
rect 684 1322 736 1332
rect 893 1322 945 1332
rect 736 1270 893 1322
rect 684 1260 736 1270
rect 893 1260 945 1270
rect -72 1236 -20 1246
rect -407 1202 -355 1212
rect -355 1184 -72 1202
rect 113 1236 165 1246
rect -20 1184 113 1202
rect 389 1236 441 1246
rect 165 1184 389 1202
rect 573 1236 625 1246
rect 441 1184 573 1202
rect 893 1202 945 1212
rect 625 1184 893 1202
rect -355 1150 893 1184
rect -407 1140 -355 1150
rect 893 1140 945 1150
rect 471 1098 529 1110
rect 471 1046 474 1098
rect 526 1046 529 1098
rect 471 1034 529 1046
rect -814 1006 -758 1016
rect -198 1006 -146 1016
rect 1534 1006 1590 1016
rect -814 954 -812 1006
rect -760 954 -198 1006
rect -146 975 1536 1006
rect -146 954 -74 975
rect -814 944 -758 954
rect -198 944 -146 954
rect -81 923 -74 954
rect -22 954 1536 975
rect 1588 954 1590 1006
rect -22 923 -14 954
rect 1534 944 1590 954
rect -81 912 -14 923
rect 548 902 615 919
rect -1052 882 -996 892
rect 548 882 555 902
rect -1052 830 -1050 882
rect -998 850 555 882
rect 607 882 615 902
rect 684 882 736 892
rect 1296 882 1352 892
rect 607 850 684 882
rect -998 830 684 850
rect 736 830 1298 882
rect 1350 830 1352 882
rect -1052 820 -996 830
rect 684 820 736 830
rect 1296 820 1352 830
rect 97 787 155 797
rect -268 785 155 787
rect -268 735 100 785
rect 97 733 100 735
rect 152 733 155 785
rect 97 721 155 733
rect 513 782 571 792
rect 513 780 806 782
rect 513 728 516 780
rect 568 728 806 780
rect 513 726 806 728
rect 513 716 571 726
rect -1174 424 -1118 434
rect -1062 424 -1006 434
rect -1174 417 -1006 424
rect -1174 365 -1172 417
rect -1120 365 -1060 417
rect -1008 365 -1006 417
rect -1174 358 -1006 365
rect -1174 348 -1118 358
rect -1062 348 -1006 358
rect 1544 424 1600 434
rect 1656 424 1712 434
rect 1544 417 1712 424
rect 1544 365 1546 417
rect 1598 365 1658 417
rect 1710 365 1712 417
rect 1544 358 1712 365
rect 1544 348 1600 358
rect 1656 348 1712 358
<< via2 >>
rect 796 1787 852 1789
rect 796 1735 798 1787
rect 798 1735 850 1787
rect 850 1735 852 1787
rect 796 1733 852 1735
rect -192 1417 -136 1473
<< metal3 >>
rect -212 1793 -116 1804
rect -212 1729 -196 1793
rect -132 1729 -116 1793
rect -212 1718 -116 1729
rect 776 1793 872 1815
rect 776 1729 792 1793
rect 856 1729 872 1793
rect -202 1473 -126 1718
rect 776 1708 872 1729
rect -202 1417 -192 1473
rect -136 1417 -126 1473
rect -202 1407 -126 1417
<< via3 >>
rect -196 1729 -132 1793
rect 792 1789 856 1793
rect 792 1733 796 1789
rect 796 1733 852 1789
rect 852 1733 856 1789
rect 792 1729 856 1733
<< metal4 >>
rect -203 1793 863 1805
rect -203 1729 -196 1793
rect -132 1729 792 1793
rect 856 1729 863 1793
rect -203 1717 863 1729
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1731262622
transform 1 0 -98 0 1 644
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1731262622
transform 1 0 360 0 1 644
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_R8XU9D  XM1
timestamp 1731262622
transform 0 1 -655 -1 0 1761
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM2
timestamp 1731262622
transform 0 -1 -655 1 0 1445
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM3
timestamp 1731262622
transform 0 1 1193 -1 0 1761
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM4
timestamp 1731262622
transform 0 1 1193 -1 0 1445
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_R8XU9D  XM5
timestamp 1731262622
transform 0 1 -655 -1 0 1129
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM6
timestamp 1731262622
transform 0 -1 -864 1 0 707
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_TGNW9T  XM7
timestamp 1731262622
transform 0 1 -864 -1 0 391
box -201 -300 201 300
use sky130_fd_pr__pfet_01v8_R8XU9D  XM8
timestamp 1731262622
transform 0 1 1193 -1 0 1129
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_TGNW9T  XM9
timestamp 1731262622
transform 0 1 1402 -1 0 707
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_TGNW9T  XM10
timestamp 1731262622
transform 0 1 1402 -1 0 391
box -201 -300 201 300
<< labels >>
flabel metal2 s -262 735 -210 787 0 FreeSans 1250 0 0 0 OUT
port 1 nsew
flabel metal2 s 750 726 806 782 0 FreeSans 1250 0 0 0 OUTN
port 2 nsew
flabel metal2 s -1118 1728 -1052 1794 0 FreeSans 1250 0 0 0 INN
port 3 nsew
flabel metal2 s -1118 1412 -1052 1478 0 FreeSans 1250 0 0 0 INP
port 4 nsew
flabel metal1 s 237 1875 336 1972 0 FreeSans 1250 0 0 0 VDD
port 5 nsew
flabel metal1 s 252 180 351 277 0 FreeSans 1250 0 0 0 VSS
port 6 nsew
<< end >>
