magic
tech sky130A
magscale 1 2
timestamp 1731262622
<< pwell >>
rect -1686 -400 1686 400
<< nmoslvt >>
rect -1500 -200 1500 200
<< ndiff >>
rect -1558 187 -1500 200
rect -1558 153 -1546 187
rect -1512 153 -1500 187
rect -1558 119 -1500 153
rect -1558 85 -1546 119
rect -1512 85 -1500 119
rect -1558 51 -1500 85
rect -1558 17 -1546 51
rect -1512 17 -1500 51
rect -1558 -17 -1500 17
rect -1558 -51 -1546 -17
rect -1512 -51 -1500 -17
rect -1558 -85 -1500 -51
rect -1558 -119 -1546 -85
rect -1512 -119 -1500 -85
rect -1558 -153 -1500 -119
rect -1558 -187 -1546 -153
rect -1512 -187 -1500 -153
rect -1558 -200 -1500 -187
rect 1500 187 1558 200
rect 1500 153 1512 187
rect 1546 153 1558 187
rect 1500 119 1558 153
rect 1500 85 1512 119
rect 1546 85 1558 119
rect 1500 51 1558 85
rect 1500 17 1512 51
rect 1546 17 1558 51
rect 1500 -17 1558 17
rect 1500 -51 1512 -17
rect 1546 -51 1558 -17
rect 1500 -85 1558 -51
rect 1500 -119 1512 -85
rect 1546 -119 1558 -85
rect 1500 -153 1558 -119
rect 1500 -187 1512 -153
rect 1546 -187 1558 -153
rect 1500 -200 1558 -187
<< ndiffc >>
rect -1546 153 -1512 187
rect -1546 85 -1512 119
rect -1546 17 -1512 51
rect -1546 -51 -1512 -17
rect -1546 -119 -1512 -85
rect -1546 -187 -1512 -153
rect 1512 153 1546 187
rect 1512 85 1546 119
rect 1512 17 1546 51
rect 1512 -51 1546 -17
rect 1512 -119 1546 -85
rect 1512 -187 1546 -153
<< psubdiff >>
rect -1660 340 -1547 374
rect -1513 340 -1479 374
rect -1445 340 -1411 374
rect -1377 340 -1343 374
rect -1309 340 -1275 374
rect -1241 340 -1207 374
rect -1173 340 -1139 374
rect -1105 340 -1071 374
rect -1037 340 -1003 374
rect -969 340 -935 374
rect -901 340 -867 374
rect -833 340 -799 374
rect -765 340 -731 374
rect -697 340 -663 374
rect -629 340 -595 374
rect -561 340 -527 374
rect -493 340 -459 374
rect -425 340 -391 374
rect -357 340 -323 374
rect -289 340 -255 374
rect -221 340 -187 374
rect -153 340 -119 374
rect -85 340 -51 374
rect -17 340 17 374
rect 51 340 85 374
rect 119 340 153 374
rect 187 340 221 374
rect 255 340 289 374
rect 323 340 357 374
rect 391 340 425 374
rect 459 340 493 374
rect 527 340 561 374
rect 595 340 629 374
rect 663 340 697 374
rect 731 340 765 374
rect 799 340 833 374
rect 867 340 901 374
rect 935 340 969 374
rect 1003 340 1037 374
rect 1071 340 1105 374
rect 1139 340 1173 374
rect 1207 340 1241 374
rect 1275 340 1309 374
rect 1343 340 1377 374
rect 1411 340 1445 374
rect 1479 340 1513 374
rect 1547 340 1660 374
rect -1660 255 -1626 340
rect -1660 187 -1626 221
rect 1626 255 1660 340
rect -1660 119 -1626 153
rect -1660 51 -1626 85
rect -1660 -17 -1626 17
rect -1660 -85 -1626 -51
rect -1660 -153 -1626 -119
rect -1660 -221 -1626 -187
rect 1626 187 1660 221
rect 1626 119 1660 153
rect 1626 51 1660 85
rect 1626 -17 1660 17
rect 1626 -85 1660 -51
rect 1626 -153 1660 -119
rect -1660 -340 -1626 -255
rect 1626 -221 1660 -187
rect 1626 -340 1660 -255
rect -1660 -374 -1547 -340
rect -1513 -374 -1479 -340
rect -1445 -374 -1411 -340
rect -1377 -374 -1343 -340
rect -1309 -374 -1275 -340
rect -1241 -374 -1207 -340
rect -1173 -374 -1139 -340
rect -1105 -374 -1071 -340
rect -1037 -374 -1003 -340
rect -969 -374 -935 -340
rect -901 -374 -867 -340
rect -833 -374 -799 -340
rect -765 -374 -731 -340
rect -697 -374 -663 -340
rect -629 -374 -595 -340
rect -561 -374 -527 -340
rect -493 -374 -459 -340
rect -425 -374 -391 -340
rect -357 -374 -323 -340
rect -289 -374 -255 -340
rect -221 -374 -187 -340
rect -153 -374 -119 -340
rect -85 -374 -51 -340
rect -17 -374 17 -340
rect 51 -374 85 -340
rect 119 -374 153 -340
rect 187 -374 221 -340
rect 255 -374 289 -340
rect 323 -374 357 -340
rect 391 -374 425 -340
rect 459 -374 493 -340
rect 527 -374 561 -340
rect 595 -374 629 -340
rect 663 -374 697 -340
rect 731 -374 765 -340
rect 799 -374 833 -340
rect 867 -374 901 -340
rect 935 -374 969 -340
rect 1003 -374 1037 -340
rect 1071 -374 1105 -340
rect 1139 -374 1173 -340
rect 1207 -374 1241 -340
rect 1275 -374 1309 -340
rect 1343 -374 1377 -340
rect 1411 -374 1445 -340
rect 1479 -374 1513 -340
rect 1547 -374 1660 -340
<< psubdiffcont >>
rect -1547 340 -1513 374
rect -1479 340 -1445 374
rect -1411 340 -1377 374
rect -1343 340 -1309 374
rect -1275 340 -1241 374
rect -1207 340 -1173 374
rect -1139 340 -1105 374
rect -1071 340 -1037 374
rect -1003 340 -969 374
rect -935 340 -901 374
rect -867 340 -833 374
rect -799 340 -765 374
rect -731 340 -697 374
rect -663 340 -629 374
rect -595 340 -561 374
rect -527 340 -493 374
rect -459 340 -425 374
rect -391 340 -357 374
rect -323 340 -289 374
rect -255 340 -221 374
rect -187 340 -153 374
rect -119 340 -85 374
rect -51 340 -17 374
rect 17 340 51 374
rect 85 340 119 374
rect 153 340 187 374
rect 221 340 255 374
rect 289 340 323 374
rect 357 340 391 374
rect 425 340 459 374
rect 493 340 527 374
rect 561 340 595 374
rect 629 340 663 374
rect 697 340 731 374
rect 765 340 799 374
rect 833 340 867 374
rect 901 340 935 374
rect 969 340 1003 374
rect 1037 340 1071 374
rect 1105 340 1139 374
rect 1173 340 1207 374
rect 1241 340 1275 374
rect 1309 340 1343 374
rect 1377 340 1411 374
rect 1445 340 1479 374
rect 1513 340 1547 374
rect -1660 221 -1626 255
rect 1626 221 1660 255
rect -1660 153 -1626 187
rect -1660 85 -1626 119
rect -1660 17 -1626 51
rect -1660 -51 -1626 -17
rect -1660 -119 -1626 -85
rect -1660 -187 -1626 -153
rect 1626 153 1660 187
rect 1626 85 1660 119
rect 1626 17 1660 51
rect 1626 -51 1660 -17
rect 1626 -119 1660 -85
rect 1626 -187 1660 -153
rect -1660 -255 -1626 -221
rect 1626 -255 1660 -221
rect -1547 -374 -1513 -340
rect -1479 -374 -1445 -340
rect -1411 -374 -1377 -340
rect -1343 -374 -1309 -340
rect -1275 -374 -1241 -340
rect -1207 -374 -1173 -340
rect -1139 -374 -1105 -340
rect -1071 -374 -1037 -340
rect -1003 -374 -969 -340
rect -935 -374 -901 -340
rect -867 -374 -833 -340
rect -799 -374 -765 -340
rect -731 -374 -697 -340
rect -663 -374 -629 -340
rect -595 -374 -561 -340
rect -527 -374 -493 -340
rect -459 -374 -425 -340
rect -391 -374 -357 -340
rect -323 -374 -289 -340
rect -255 -374 -221 -340
rect -187 -374 -153 -340
rect -119 -374 -85 -340
rect -51 -374 -17 -340
rect 17 -374 51 -340
rect 85 -374 119 -340
rect 153 -374 187 -340
rect 221 -374 255 -340
rect 289 -374 323 -340
rect 357 -374 391 -340
rect 425 -374 459 -340
rect 493 -374 527 -340
rect 561 -374 595 -340
rect 629 -374 663 -340
rect 697 -374 731 -340
rect 765 -374 799 -340
rect 833 -374 867 -340
rect 901 -374 935 -340
rect 969 -374 1003 -340
rect 1037 -374 1071 -340
rect 1105 -374 1139 -340
rect 1173 -374 1207 -340
rect 1241 -374 1275 -340
rect 1309 -374 1343 -340
rect 1377 -374 1411 -340
rect 1445 -374 1479 -340
rect 1513 -374 1547 -340
<< poly >>
rect -1500 272 1500 288
rect -1500 238 -1479 272
rect -1445 238 -1411 272
rect -1377 238 -1343 272
rect -1309 238 -1275 272
rect -1241 238 -1207 272
rect -1173 238 -1139 272
rect -1105 238 -1071 272
rect -1037 238 -1003 272
rect -969 238 -935 272
rect -901 238 -867 272
rect -833 238 -799 272
rect -765 238 -731 272
rect -697 238 -663 272
rect -629 238 -595 272
rect -561 238 -527 272
rect -493 238 -459 272
rect -425 238 -391 272
rect -357 238 -323 272
rect -289 238 -255 272
rect -221 238 -187 272
rect -153 238 -119 272
rect -85 238 -51 272
rect -17 238 17 272
rect 51 238 85 272
rect 119 238 153 272
rect 187 238 221 272
rect 255 238 289 272
rect 323 238 357 272
rect 391 238 425 272
rect 459 238 493 272
rect 527 238 561 272
rect 595 238 629 272
rect 663 238 697 272
rect 731 238 765 272
rect 799 238 833 272
rect 867 238 901 272
rect 935 238 969 272
rect 1003 238 1037 272
rect 1071 238 1105 272
rect 1139 238 1173 272
rect 1207 238 1241 272
rect 1275 238 1309 272
rect 1343 238 1377 272
rect 1411 238 1445 272
rect 1479 238 1500 272
rect -1500 200 1500 238
rect -1500 -238 1500 -200
rect -1500 -272 -1479 -238
rect -1445 -272 -1411 -238
rect -1377 -272 -1343 -238
rect -1309 -272 -1275 -238
rect -1241 -272 -1207 -238
rect -1173 -272 -1139 -238
rect -1105 -272 -1071 -238
rect -1037 -272 -1003 -238
rect -969 -272 -935 -238
rect -901 -272 -867 -238
rect -833 -272 -799 -238
rect -765 -272 -731 -238
rect -697 -272 -663 -238
rect -629 -272 -595 -238
rect -561 -272 -527 -238
rect -493 -272 -459 -238
rect -425 -272 -391 -238
rect -357 -272 -323 -238
rect -289 -272 -255 -238
rect -221 -272 -187 -238
rect -153 -272 -119 -238
rect -85 -272 -51 -238
rect -17 -272 17 -238
rect 51 -272 85 -238
rect 119 -272 153 -238
rect 187 -272 221 -238
rect 255 -272 289 -238
rect 323 -272 357 -238
rect 391 -272 425 -238
rect 459 -272 493 -238
rect 527 -272 561 -238
rect 595 -272 629 -238
rect 663 -272 697 -238
rect 731 -272 765 -238
rect 799 -272 833 -238
rect 867 -272 901 -238
rect 935 -272 969 -238
rect 1003 -272 1037 -238
rect 1071 -272 1105 -238
rect 1139 -272 1173 -238
rect 1207 -272 1241 -238
rect 1275 -272 1309 -238
rect 1343 -272 1377 -238
rect 1411 -272 1445 -238
rect 1479 -272 1500 -238
rect -1500 -288 1500 -272
<< polycont >>
rect -1479 238 -1445 272
rect -1411 238 -1377 272
rect -1343 238 -1309 272
rect -1275 238 -1241 272
rect -1207 238 -1173 272
rect -1139 238 -1105 272
rect -1071 238 -1037 272
rect -1003 238 -969 272
rect -935 238 -901 272
rect -867 238 -833 272
rect -799 238 -765 272
rect -731 238 -697 272
rect -663 238 -629 272
rect -595 238 -561 272
rect -527 238 -493 272
rect -459 238 -425 272
rect -391 238 -357 272
rect -323 238 -289 272
rect -255 238 -221 272
rect -187 238 -153 272
rect -119 238 -85 272
rect -51 238 -17 272
rect 17 238 51 272
rect 85 238 119 272
rect 153 238 187 272
rect 221 238 255 272
rect 289 238 323 272
rect 357 238 391 272
rect 425 238 459 272
rect 493 238 527 272
rect 561 238 595 272
rect 629 238 663 272
rect 697 238 731 272
rect 765 238 799 272
rect 833 238 867 272
rect 901 238 935 272
rect 969 238 1003 272
rect 1037 238 1071 272
rect 1105 238 1139 272
rect 1173 238 1207 272
rect 1241 238 1275 272
rect 1309 238 1343 272
rect 1377 238 1411 272
rect 1445 238 1479 272
rect -1479 -272 -1445 -238
rect -1411 -272 -1377 -238
rect -1343 -272 -1309 -238
rect -1275 -272 -1241 -238
rect -1207 -272 -1173 -238
rect -1139 -272 -1105 -238
rect -1071 -272 -1037 -238
rect -1003 -272 -969 -238
rect -935 -272 -901 -238
rect -867 -272 -833 -238
rect -799 -272 -765 -238
rect -731 -272 -697 -238
rect -663 -272 -629 -238
rect -595 -272 -561 -238
rect -527 -272 -493 -238
rect -459 -272 -425 -238
rect -391 -272 -357 -238
rect -323 -272 -289 -238
rect -255 -272 -221 -238
rect -187 -272 -153 -238
rect -119 -272 -85 -238
rect -51 -272 -17 -238
rect 17 -272 51 -238
rect 85 -272 119 -238
rect 153 -272 187 -238
rect 221 -272 255 -238
rect 289 -272 323 -238
rect 357 -272 391 -238
rect 425 -272 459 -238
rect 493 -272 527 -238
rect 561 -272 595 -238
rect 629 -272 663 -238
rect 697 -272 731 -238
rect 765 -272 799 -238
rect 833 -272 867 -238
rect 901 -272 935 -238
rect 969 -272 1003 -238
rect 1037 -272 1071 -238
rect 1105 -272 1139 -238
rect 1173 -272 1207 -238
rect 1241 -272 1275 -238
rect 1309 -272 1343 -238
rect 1377 -272 1411 -238
rect 1445 -272 1479 -238
<< locali >>
rect -1660 340 -1547 374
rect -1513 340 -1479 374
rect -1445 340 -1411 374
rect -1377 340 -1343 374
rect -1309 340 -1275 374
rect -1241 340 -1207 374
rect -1173 340 -1139 374
rect -1105 340 -1071 374
rect -1037 340 -1003 374
rect -969 340 -935 374
rect -901 340 -867 374
rect -833 340 -799 374
rect -765 340 -731 374
rect -697 340 -663 374
rect -629 340 -595 374
rect -561 340 -527 374
rect -493 340 -459 374
rect -425 340 -391 374
rect -357 340 -323 374
rect -289 340 -255 374
rect -221 340 -187 374
rect -153 340 -119 374
rect -85 340 -51 374
rect -17 340 17 374
rect 51 340 85 374
rect 119 340 153 374
rect 187 340 221 374
rect 255 340 289 374
rect 323 340 357 374
rect 391 340 425 374
rect 459 340 493 374
rect 527 340 561 374
rect 595 340 629 374
rect 663 340 697 374
rect 731 340 765 374
rect 799 340 833 374
rect 867 340 901 374
rect 935 340 969 374
rect 1003 340 1037 374
rect 1071 340 1105 374
rect 1139 340 1173 374
rect 1207 340 1241 374
rect 1275 340 1309 374
rect 1343 340 1377 374
rect 1411 340 1445 374
rect 1479 340 1513 374
rect 1547 340 1660 374
rect -1660 255 -1626 340
rect -1500 238 -1479 272
rect -1423 238 -1411 272
rect -1351 238 -1343 272
rect -1279 238 -1275 272
rect -1173 238 -1169 272
rect -1105 238 -1097 272
rect -1037 238 -1025 272
rect -969 238 -953 272
rect -901 238 -881 272
rect -833 238 -809 272
rect -765 238 -737 272
rect -697 238 -665 272
rect -629 238 -595 272
rect -559 238 -527 272
rect -487 238 -459 272
rect -415 238 -391 272
rect -343 238 -323 272
rect -271 238 -255 272
rect -199 238 -187 272
rect -127 238 -119 272
rect -55 238 -51 272
rect 51 238 55 272
rect 119 238 127 272
rect 187 238 199 272
rect 255 238 271 272
rect 323 238 343 272
rect 391 238 415 272
rect 459 238 487 272
rect 527 238 559 272
rect 595 238 629 272
rect 665 238 697 272
rect 737 238 765 272
rect 809 238 833 272
rect 881 238 901 272
rect 953 238 969 272
rect 1025 238 1037 272
rect 1097 238 1105 272
rect 1169 238 1173 272
rect 1275 238 1279 272
rect 1343 238 1351 272
rect 1411 238 1423 272
rect 1479 238 1500 272
rect 1626 255 1660 340
rect -1660 187 -1626 221
rect -1660 119 -1626 153
rect -1660 51 -1626 85
rect -1660 -17 -1626 17
rect -1660 -85 -1626 -51
rect -1660 -153 -1626 -119
rect -1660 -221 -1626 -187
rect -1546 187 -1512 204
rect -1546 119 -1512 127
rect -1546 51 -1512 55
rect -1546 -55 -1512 -51
rect -1546 -127 -1512 -119
rect -1546 -204 -1512 -187
rect 1512 187 1546 204
rect 1512 119 1546 127
rect 1512 51 1546 55
rect 1512 -55 1546 -51
rect 1512 -127 1546 -119
rect 1512 -204 1546 -187
rect 1626 187 1660 221
rect 1626 119 1660 153
rect 1626 51 1660 85
rect 1626 -17 1660 17
rect 1626 -85 1660 -51
rect 1626 -153 1660 -119
rect 1626 -221 1660 -187
rect -1660 -340 -1626 -255
rect -1500 -272 -1479 -238
rect -1423 -272 -1411 -238
rect -1351 -272 -1343 -238
rect -1279 -272 -1275 -238
rect -1173 -272 -1169 -238
rect -1105 -272 -1097 -238
rect -1037 -272 -1025 -238
rect -969 -272 -953 -238
rect -901 -272 -881 -238
rect -833 -272 -809 -238
rect -765 -272 -737 -238
rect -697 -272 -665 -238
rect -629 -272 -595 -238
rect -559 -272 -527 -238
rect -487 -272 -459 -238
rect -415 -272 -391 -238
rect -343 -272 -323 -238
rect -271 -272 -255 -238
rect -199 -272 -187 -238
rect -127 -272 -119 -238
rect -55 -272 -51 -238
rect 51 -272 55 -238
rect 119 -272 127 -238
rect 187 -272 199 -238
rect 255 -272 271 -238
rect 323 -272 343 -238
rect 391 -272 415 -238
rect 459 -272 487 -238
rect 527 -272 559 -238
rect 595 -272 629 -238
rect 665 -272 697 -238
rect 737 -272 765 -238
rect 809 -272 833 -238
rect 881 -272 901 -238
rect 953 -272 969 -238
rect 1025 -272 1037 -238
rect 1097 -272 1105 -238
rect 1169 -272 1173 -238
rect 1275 -272 1279 -238
rect 1343 -272 1351 -238
rect 1411 -272 1423 -238
rect 1479 -272 1500 -238
rect 1626 -340 1660 -255
rect -1660 -374 -1547 -340
rect -1513 -374 -1479 -340
rect -1445 -374 -1411 -340
rect -1377 -374 -1343 -340
rect -1309 -374 -1275 -340
rect -1241 -374 -1207 -340
rect -1173 -374 -1139 -340
rect -1105 -374 -1071 -340
rect -1037 -374 -1003 -340
rect -969 -374 -935 -340
rect -901 -374 -867 -340
rect -833 -374 -799 -340
rect -765 -374 -731 -340
rect -697 -374 -663 -340
rect -629 -374 -595 -340
rect -561 -374 -527 -340
rect -493 -374 -459 -340
rect -425 -374 -391 -340
rect -357 -374 -323 -340
rect -289 -374 -255 -340
rect -221 -374 -187 -340
rect -153 -374 -119 -340
rect -85 -374 -51 -340
rect -17 -374 17 -340
rect 51 -374 85 -340
rect 119 -374 153 -340
rect 187 -374 221 -340
rect 255 -374 289 -340
rect 323 -374 357 -340
rect 391 -374 425 -340
rect 459 -374 493 -340
rect 527 -374 561 -340
rect 595 -374 629 -340
rect 663 -374 697 -340
rect 731 -374 765 -340
rect 799 -374 833 -340
rect 867 -374 901 -340
rect 935 -374 969 -340
rect 1003 -374 1037 -340
rect 1071 -374 1105 -340
rect 1139 -374 1173 -340
rect 1207 -374 1241 -340
rect 1275 -374 1309 -340
rect 1343 -374 1377 -340
rect 1411 -374 1445 -340
rect 1479 -374 1513 -340
rect 1547 -374 1660 -340
<< viali >>
rect -1457 238 -1445 272
rect -1445 238 -1423 272
rect -1385 238 -1377 272
rect -1377 238 -1351 272
rect -1313 238 -1309 272
rect -1309 238 -1279 272
rect -1241 238 -1207 272
rect -1169 238 -1139 272
rect -1139 238 -1135 272
rect -1097 238 -1071 272
rect -1071 238 -1063 272
rect -1025 238 -1003 272
rect -1003 238 -991 272
rect -953 238 -935 272
rect -935 238 -919 272
rect -881 238 -867 272
rect -867 238 -847 272
rect -809 238 -799 272
rect -799 238 -775 272
rect -737 238 -731 272
rect -731 238 -703 272
rect -665 238 -663 272
rect -663 238 -631 272
rect -593 238 -561 272
rect -561 238 -559 272
rect -521 238 -493 272
rect -493 238 -487 272
rect -449 238 -425 272
rect -425 238 -415 272
rect -377 238 -357 272
rect -357 238 -343 272
rect -305 238 -289 272
rect -289 238 -271 272
rect -233 238 -221 272
rect -221 238 -199 272
rect -161 238 -153 272
rect -153 238 -127 272
rect -89 238 -85 272
rect -85 238 -55 272
rect -17 238 17 272
rect 55 238 85 272
rect 85 238 89 272
rect 127 238 153 272
rect 153 238 161 272
rect 199 238 221 272
rect 221 238 233 272
rect 271 238 289 272
rect 289 238 305 272
rect 343 238 357 272
rect 357 238 377 272
rect 415 238 425 272
rect 425 238 449 272
rect 487 238 493 272
rect 493 238 521 272
rect 559 238 561 272
rect 561 238 593 272
rect 631 238 663 272
rect 663 238 665 272
rect 703 238 731 272
rect 731 238 737 272
rect 775 238 799 272
rect 799 238 809 272
rect 847 238 867 272
rect 867 238 881 272
rect 919 238 935 272
rect 935 238 953 272
rect 991 238 1003 272
rect 1003 238 1025 272
rect 1063 238 1071 272
rect 1071 238 1097 272
rect 1135 238 1139 272
rect 1139 238 1169 272
rect 1207 238 1241 272
rect 1279 238 1309 272
rect 1309 238 1313 272
rect 1351 238 1377 272
rect 1377 238 1385 272
rect 1423 238 1445 272
rect 1445 238 1457 272
rect -1546 153 -1512 161
rect -1546 127 -1512 153
rect -1546 85 -1512 89
rect -1546 55 -1512 85
rect -1546 -17 -1512 17
rect -1546 -85 -1512 -55
rect -1546 -89 -1512 -85
rect -1546 -153 -1512 -127
rect -1546 -161 -1512 -153
rect 1512 153 1546 161
rect 1512 127 1546 153
rect 1512 85 1546 89
rect 1512 55 1546 85
rect 1512 -17 1546 17
rect 1512 -85 1546 -55
rect 1512 -89 1546 -85
rect 1512 -153 1546 -127
rect 1512 -161 1546 -153
rect -1457 -272 -1445 -238
rect -1445 -272 -1423 -238
rect -1385 -272 -1377 -238
rect -1377 -272 -1351 -238
rect -1313 -272 -1309 -238
rect -1309 -272 -1279 -238
rect -1241 -272 -1207 -238
rect -1169 -272 -1139 -238
rect -1139 -272 -1135 -238
rect -1097 -272 -1071 -238
rect -1071 -272 -1063 -238
rect -1025 -272 -1003 -238
rect -1003 -272 -991 -238
rect -953 -272 -935 -238
rect -935 -272 -919 -238
rect -881 -272 -867 -238
rect -867 -272 -847 -238
rect -809 -272 -799 -238
rect -799 -272 -775 -238
rect -737 -272 -731 -238
rect -731 -272 -703 -238
rect -665 -272 -663 -238
rect -663 -272 -631 -238
rect -593 -272 -561 -238
rect -561 -272 -559 -238
rect -521 -272 -493 -238
rect -493 -272 -487 -238
rect -449 -272 -425 -238
rect -425 -272 -415 -238
rect -377 -272 -357 -238
rect -357 -272 -343 -238
rect -305 -272 -289 -238
rect -289 -272 -271 -238
rect -233 -272 -221 -238
rect -221 -272 -199 -238
rect -161 -272 -153 -238
rect -153 -272 -127 -238
rect -89 -272 -85 -238
rect -85 -272 -55 -238
rect -17 -272 17 -238
rect 55 -272 85 -238
rect 85 -272 89 -238
rect 127 -272 153 -238
rect 153 -272 161 -238
rect 199 -272 221 -238
rect 221 -272 233 -238
rect 271 -272 289 -238
rect 289 -272 305 -238
rect 343 -272 357 -238
rect 357 -272 377 -238
rect 415 -272 425 -238
rect 425 -272 449 -238
rect 487 -272 493 -238
rect 493 -272 521 -238
rect 559 -272 561 -238
rect 561 -272 593 -238
rect 631 -272 663 -238
rect 663 -272 665 -238
rect 703 -272 731 -238
rect 731 -272 737 -238
rect 775 -272 799 -238
rect 799 -272 809 -238
rect 847 -272 867 -238
rect 867 -272 881 -238
rect 919 -272 935 -238
rect 935 -272 953 -238
rect 991 -272 1003 -238
rect 1003 -272 1025 -238
rect 1063 -272 1071 -238
rect 1071 -272 1097 -238
rect 1135 -272 1139 -238
rect 1139 -272 1169 -238
rect 1207 -272 1241 -238
rect 1279 -272 1309 -238
rect 1309 -272 1313 -238
rect 1351 -272 1377 -238
rect 1377 -272 1385 -238
rect 1423 -272 1445 -238
rect 1445 -272 1457 -238
<< metal1 >>
rect -1496 272 1496 278
rect -1496 238 -1457 272
rect -1423 238 -1385 272
rect -1351 238 -1313 272
rect -1279 238 -1241 272
rect -1207 238 -1169 272
rect -1135 238 -1097 272
rect -1063 238 -1025 272
rect -991 238 -953 272
rect -919 238 -881 272
rect -847 238 -809 272
rect -775 238 -737 272
rect -703 238 -665 272
rect -631 238 -593 272
rect -559 238 -521 272
rect -487 238 -449 272
rect -415 238 -377 272
rect -343 238 -305 272
rect -271 238 -233 272
rect -199 238 -161 272
rect -127 238 -89 272
rect -55 238 -17 272
rect 17 238 55 272
rect 89 238 127 272
rect 161 238 199 272
rect 233 238 271 272
rect 305 238 343 272
rect 377 238 415 272
rect 449 238 487 272
rect 521 238 559 272
rect 593 238 631 272
rect 665 238 703 272
rect 737 238 775 272
rect 809 238 847 272
rect 881 238 919 272
rect 953 238 991 272
rect 1025 238 1063 272
rect 1097 238 1135 272
rect 1169 238 1207 272
rect 1241 238 1279 272
rect 1313 238 1351 272
rect 1385 238 1423 272
rect 1457 238 1496 272
rect -1496 232 1496 238
rect -1552 161 -1506 200
rect -1552 127 -1546 161
rect -1512 127 -1506 161
rect -1552 89 -1506 127
rect -1552 55 -1546 89
rect -1512 55 -1506 89
rect -1552 17 -1506 55
rect -1552 -17 -1546 17
rect -1512 -17 -1506 17
rect -1552 -55 -1506 -17
rect -1552 -89 -1546 -55
rect -1512 -89 -1506 -55
rect -1552 -127 -1506 -89
rect -1552 -161 -1546 -127
rect -1512 -161 -1506 -127
rect -1552 -200 -1506 -161
rect 1506 161 1552 200
rect 1506 127 1512 161
rect 1546 127 1552 161
rect 1506 89 1552 127
rect 1506 55 1512 89
rect 1546 55 1552 89
rect 1506 17 1552 55
rect 1506 -17 1512 17
rect 1546 -17 1552 17
rect 1506 -55 1552 -17
rect 1506 -89 1512 -55
rect 1546 -89 1552 -55
rect 1506 -127 1552 -89
rect 1506 -161 1512 -127
rect 1546 -161 1552 -127
rect 1506 -200 1552 -161
rect -1496 -238 1496 -232
rect -1496 -272 -1457 -238
rect -1423 -272 -1385 -238
rect -1351 -272 -1313 -238
rect -1279 -272 -1241 -238
rect -1207 -272 -1169 -238
rect -1135 -272 -1097 -238
rect -1063 -272 -1025 -238
rect -991 -272 -953 -238
rect -919 -272 -881 -238
rect -847 -272 -809 -238
rect -775 -272 -737 -238
rect -703 -272 -665 -238
rect -631 -272 -593 -238
rect -559 -272 -521 -238
rect -487 -272 -449 -238
rect -415 -272 -377 -238
rect -343 -272 -305 -238
rect -271 -272 -233 -238
rect -199 -272 -161 -238
rect -127 -272 -89 -238
rect -55 -272 -17 -238
rect 17 -272 55 -238
rect 89 -272 127 -238
rect 161 -272 199 -238
rect 233 -272 271 -238
rect 305 -272 343 -238
rect 377 -272 415 -238
rect 449 -272 487 -238
rect 521 -272 559 -238
rect 593 -272 631 -238
rect 665 -272 703 -238
rect 737 -272 775 -238
rect 809 -272 847 -238
rect 881 -272 919 -238
rect 953 -272 991 -238
rect 1025 -272 1063 -238
rect 1097 -272 1135 -238
rect 1169 -272 1207 -238
rect 1241 -272 1279 -238
rect 1313 -272 1351 -238
rect 1385 -272 1423 -238
rect 1457 -272 1496 -238
rect -1496 -278 1496 -272
<< properties >>
string FIXED_BBOX -1642 -356 1642 356
<< end >>
