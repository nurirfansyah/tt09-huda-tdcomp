magic
tech sky130A
magscale 1 2
timestamp 1731262622
<< nwell >>
rect 24654 16815 26560 16831
rect 24267 15777 26560 16815
rect 25434 14984 26000 15777
<< metal1 >>
rect 22638 17700 23058 17714
rect 22638 17328 22662 17700
rect 23034 17328 23058 17700
rect 22638 17314 23058 17328
<< via1 >>
rect 22662 17328 23034 17700
<< metal2 >>
rect 26209 17818 26308 17849
rect 25135 17768 25234 17799
rect 22648 17702 23048 17724
rect 22648 17326 22660 17702
rect 23036 17326 23048 17702
rect 25135 17712 25156 17768
rect 25212 17712 25234 17768
rect 26209 17762 26230 17818
rect 26286 17762 26308 17818
rect 26209 17732 26308 17762
rect 25135 17682 25234 17712
rect 22648 17304 23048 17326
rect 21970 15990 22370 16012
rect 21970 15614 21982 15990
rect 22358 15614 22370 15990
rect 21970 15592 22370 15614
rect 22090 2300 22185 15592
rect 27660 4114 27782 4156
rect 27660 4058 27693 4114
rect 27749 4058 27782 4114
rect 27660 4016 27782 4058
rect 25510 3777 25612 3805
rect 25510 3721 25533 3777
rect 25589 3721 25612 3777
rect 25510 3694 25612 3721
rect 25672 2300 25767 3821
rect 25826 3777 25928 3805
rect 25826 3721 25849 3777
rect 25905 3721 25928 3777
rect 25826 3694 25928 3721
rect 22090 2205 25767 2300
<< via2 >>
rect 22660 17700 23036 17702
rect 22660 17328 22662 17700
rect 22662 17328 23034 17700
rect 23034 17328 23036 17700
rect 22660 17326 23036 17328
rect 25156 17712 25212 17768
rect 26230 17762 26286 17818
rect 21982 15614 22358 15990
rect 27693 4058 27749 4114
rect 25533 3721 25589 3777
rect 25849 3721 25905 3777
<< metal3 >>
rect 26199 17822 26318 17844
rect 25125 17772 25244 17794
rect 22638 17706 23058 17719
rect 22638 17322 22656 17706
rect 23040 17322 23058 17706
rect 25125 17708 25152 17772
rect 25216 17708 25244 17772
rect 26199 17758 26226 17822
rect 26290 17758 26318 17822
rect 26199 17737 26318 17758
rect 25125 17687 25244 17708
rect 22638 17309 23058 17322
rect 21960 15994 22380 16007
rect 21960 15610 21978 15994
rect 22362 15610 22380 15994
rect 21960 15597 22380 15610
rect 27650 4118 27792 4151
rect 27650 4054 27689 4118
rect 27753 4054 27792 4118
rect 27650 4021 27792 4054
rect 25500 3781 25622 3800
rect 25500 3717 25529 3781
rect 25593 3717 25622 3781
rect 25500 3699 25622 3717
rect 25816 3781 25938 3800
rect 25816 3717 25845 3781
rect 25909 3717 25938 3781
rect 25816 3699 25938 3717
<< via3 >>
rect 22656 17702 23040 17706
rect 22656 17326 22660 17702
rect 22660 17326 23036 17702
rect 23036 17326 23040 17702
rect 22656 17322 23040 17326
rect 25152 17768 25216 17772
rect 25152 17712 25156 17768
rect 25156 17712 25212 17768
rect 25212 17712 25216 17768
rect 25152 17708 25216 17712
rect 26226 17818 26290 17822
rect 26226 17762 26230 17818
rect 26230 17762 26286 17818
rect 26286 17762 26290 17818
rect 26226 17758 26290 17762
rect 21978 15990 22362 15994
rect 21978 15614 21982 15990
rect 21982 15614 22358 15990
rect 22358 15614 22362 15990
rect 21978 15610 22362 15614
rect 27689 4114 27753 4118
rect 27689 4058 27693 4114
rect 27693 4058 27749 4114
rect 27749 4058 27753 4114
rect 27689 4054 27753 4058
rect 25529 3777 25593 3781
rect 25529 3721 25533 3777
rect 25533 3721 25589 3777
rect 25589 3721 25593 3777
rect 25529 3717 25593 3721
rect 25845 3777 25909 3781
rect 25845 3721 25849 3777
rect 25849 3721 25905 3777
rect 25905 3721 25909 3777
rect 25845 3717 25909 3721
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 200 16002 600 44152
rect 800 17714 1200 44152
rect 18278 18373 18338 45152
rect 18830 18813 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 18830 18753 26289 18813
rect 18278 18313 25214 18373
rect 25154 17790 25214 18313
rect 26229 17840 26289 18753
rect 26208 17822 26309 17840
rect 25134 17772 25235 17790
rect 22647 17714 23049 17715
rect 800 17706 23049 17714
rect 800 17322 22656 17706
rect 23040 17322 23049 17706
rect 25134 17708 25152 17772
rect 25216 17708 25235 17772
rect 26208 17758 26226 17822
rect 26290 17758 26309 17822
rect 26208 17741 26309 17758
rect 25134 17691 25235 17708
rect 800 17314 23049 17322
rect 800 16002 1200 17314
rect 22647 17313 23049 17314
rect 21969 16002 22371 16003
rect 200 15994 22371 16002
rect 200 15610 21978 15994
rect 22362 15610 22371 15994
rect 200 15602 22371 15610
rect 200 1000 600 15602
rect 800 1000 1200 15602
rect 21969 15601 22371 15602
rect 27659 4118 27783 4147
rect 27659 4054 27689 4118
rect 27753 4105 27783 4118
rect 28766 4105 28826 45152
rect 29318 44952 29378 45152
rect 27753 4054 28826 4105
rect 27659 4045 28826 4054
rect 27659 4025 27783 4045
rect 25470 3781 25650 3854
rect 25470 3717 25529 3781
rect 25593 3717 25650 3781
rect 25470 2706 25650 3717
rect 25789 3781 25969 3851
rect 25789 3717 25845 3781
rect 25909 3717 25969 3781
rect 25789 3082 25969 3717
rect 25789 2902 30542 3082
rect 25470 2526 26678 2706
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 2526
rect 30362 0 30542 2902
use tdc  tdc_0
timestamp 1731262622
transform 0 -1 24988 1 0 8540
box -4836 -3737 9311 2274
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 750 90 0 0 clk
port 1 nsew
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 750 90 0 0 ena
port 2 nsew
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 750 90 0 0 rst_n
port 3 nsew
flabel metal4 s 30362 0 30542 200 0 FreeSans 1500 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26498 0 26678 200 0 FreeSans 1500 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 22634 0 22814 200 0 FreeSans 1500 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 18770 0 18950 200 0 FreeSans 1500 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 14906 0 15086 200 0 FreeSans 1500 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 11042 0 11222 200 0 FreeSans 1500 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 7178 0 7358 200 0 FreeSans 1500 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 3314 0 3494 200 0 FreeSans 1500 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 750 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 750 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 750 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 750 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 750 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 750 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 750 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 750 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 750 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 750 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 750 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 750 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 750 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 750 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 750 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 750 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 750 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 750 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 750 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 750 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 750 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 750 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 750 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 750 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 750 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 750 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 750 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 750 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 750 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 750 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 750 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 750 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 750 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 750 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 750 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 750 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 750 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 750 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 750 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 750 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 200 1000 600 44152 1 FreeSans 625 0 0 0 VDPWR
port 52 nsew
flabel metal4 s 800 1000 1200 44152 1 FreeSans 625 0 0 0 VGND
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
